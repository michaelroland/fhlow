--------------------------------------------------------------------------------
-- This file is part of fhlow (fast handling of a lot of work), a working
-- environment that speeds up the development of and structures FPGA design
-- projects.
-- 
-- Copyright (c) 2011-2016 Michael Roland <michael.roland@fh-hagenberg.at>
-- 
-- This program is free software: you can redistribute it and/or modify
-- it under the terms of the GNU General Public License as published by
-- the Free Software Foundation, either version 3 of the License, or
-- (at your option) any later version.
-- 
-- This program is distributed in the hope that it will be useful,
-- but WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
-- GNU General Public License for more details.
-- 
-- You should have received a copy of the GNU General Public License
-- along with this program.  If not, see <http://www.gnu.org/licenses/>.
--------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library example_library;
use example_library.ExamplePackage.all;

entity Example1 is
  
  port (
    iClk         : in std_ulogic;
    inResetAsync : in std_ulogic;

    oSEG0        : out std_ulogic_vector(6 downto 0);
    oSEG1        : out std_ulogic_vector(6 downto 0);
    oSEG2        : out std_ulogic_vector(6 downto 0);
    oSEG3        : out std_ulogic_vector(6 downto 0);
    oSEG4        : out std_ulogic_vector(6 downto 0);
    oSEG5        : out std_ulogic_vector(6 downto 0));

end Example1;
